/*module magic(clk, LED[9:0])

	//nightrider rules!

endmodule
*/