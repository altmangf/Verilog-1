//scratch

/*
module Project1_top(SW, KEY, HEX0, HEX1, LED);

	input [9:0]SW;
	input [1:0]Key;
	output[8:0]HEX0;
	output[9:0]HEX1;
	output[9:0]LED;
	
	wire[7:0] hexDisplay;
	
	*/