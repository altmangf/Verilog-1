/*
Gabriel Altman
ECEN 2350 Digital Logic
March, 2018
*/

/*module magic(clk, LED[9:0])

	//nightrider rules!

endmodule
*/