/*
module logicalEqual(x, y, boolean)
	output reg boolean;
	
	always @(x,y)
		begin
			if (x == y) boolean=1;
			else boolean=0;
endmodule
*/		