/*module max(x, y, xMax, yMax)
	input [3:0]x, [3:0]y;
	output reg xMax, yMax;
	
	//This module will probably use a Four-bit Magnitude Comparator
	
endmodule
*/