/*
Gabriel Altman
ECEN 2350 Digital Logic
March, 2018
*/


/*module Subtract(carryin, X, Y, S, carryout);
	parameter n=4;
	
	//subtraction code goes here.
	//n-bit Full Subtractor with parameters, For Loop, Integer statement
		
endmodule
*/