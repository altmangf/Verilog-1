/*module greater(x, y, boolean)
	input [3:0]x, [3:0]y;
	output reg boolean;
	
	always @(x,y)
		begin
			if (x > y) boolean=1;
			else boolean=0;
endmodule*/